
`define SRAM 0
`define SRAM_BITS  24
`define SRAM_BASE  8'h80

`define UART 1
`define UART_BITS  16
`define UART_BASE  16'hA000

`define ACCEL 2
`define ACCEL_BITS 16
`define ACCEL_BASE 16'h7000

`define TIMER 3
`define TIMER_BITS 16
`define TIMER_BASE 16'h6000
