module foo;

endmodule
